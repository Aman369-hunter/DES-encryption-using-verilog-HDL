`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.02.2026 17:16:29
// Design Name: 
// Module Name: sbox6
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sbox6(
    input [5:0] in,
    output reg [3:0] out
    );
    wire [1:0] row;
    wire [3:0] column;
    
    //assign 5th and 0th bit to the row
    //assign 4 to 1 bit the column
    assign row= {in[5], in[0]};
    assign column= in[4:1];
    
    always @(*) begin
    case({row,column})
    
6'b000000: out=4'd12; 6'b000001: out=4'd1;  6'b000010: out=4'd10; 6'b000011: out=4'd15;
6'b000100: out=4'd9;  6'b000101: out=4'd2;  6'b000110: out=4'd6;  6'b000111: out=4'd8;
6'b001000: out=4'd0;  6'b001001: out=4'd13; 6'b001010: out=4'd3;  6'b001011: out=4'd4;
6'b001100: out=4'd14; 6'b001101: out=4'd7;  6'b001110: out=4'd5;  6'b001111: out=4'd11;

6'b010000: out=4'd10; 6'b010001: out=4'd15; 6'b010010: out=4'd4;  6'b010011: out=4'd2;
6'b010100: out=4'd7;  6'b010101: out=4'd12; 6'b010110: out=4'd9;  6'b010111: out=4'd5;
6'b011000: out=4'd6;  6'b011001: out=4'd1;  6'b011010: out=4'd13; 6'b011011: out=4'd14;
6'b011100: out=4'd0;  6'b011101: out=4'd11; 6'b011110: out=4'd3;  6'b011111: out=4'd8;

6'b100000: out=4'd9;  6'b100001: out=4'd14; 6'b100010: out=4'd15; 6'b100011: out=4'd5;
6'b100100: out=4'd2;  6'b100101: out=4'd8;  6'b100110: out=4'd12; 6'b100111: out=4'd3;
6'b101000: out=4'd7;  6'b101001: out=4'd0;  6'b101010: out=4'd4;  6'b101011: out=4'd10;
6'b101100: out=4'd1;  6'b101101: out=4'd13; 6'b101110: out=4'd11; 6'b101111: out=4'd6;

6'b110000: out=4'd4;  6'b110001: out=4'd3;  6'b110010: out=4'd2;  6'b110011: out=4'd12;
6'b110100: out=4'd9;  6'b110101: out=4'd5;  6'b110110: out=4'd15; 6'b110111: out=4'd10;
6'b111000: out=4'd11; 6'b111001: out=4'd14; 6'b111010: out=4'd1;  6'b111011: out=4'd7;
6'b111100: out=4'd6;  6'b111101: out=4'd0;  6'b111110: out=4'd8;  6'b111111: out=4'd13;
    endcase
   end
endmodule
